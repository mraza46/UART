package my_package;

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "seq_item.sv"
  `include "seq.sv"
  `include "sequencer.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "agent.sv"
  `include "scoreboard.sv"
  `include "env.sv"
  `include "test.sv"

endpackage

